EX2                 ;标题
VS 1 0 10           ;电源 10V，连接在节点 1 和节点 0
R1 1 2 20           ;电阻 R1，20 欧姆,连接在节点 1 和节点 2
R2 2 0 20           ;电阻 R2，20 欧姆,连接在节点 2 和节点 0
R3 3 0 4000         ;电阻 R3，4k 欧姆,连接在节点 3 和节点 0
C1 3 0 0.0000005     ;电容 C，0.5 微法连接在节点 3 和节点 0
L1 2 3 0.2           ;电感 L，0.2 H,连接在节点 2 和节点 3
.TRAN 0.1M 30M UIC  ;瞬态分析,打印时间间隔 0.1ms，终止时间 30ms，使用初始化条件
.END                ;结束